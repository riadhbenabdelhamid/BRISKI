// Lookup table generated from CSV
`ifndef MMCM_LOOKUP_PARAMS_SVH
`define MMCM_LOOKUP_PARAMS_SVH

localparam int desired_freqs[638] = {
100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318, 319, 320, 321, 322, 323, 324, 325, 326, 327, 328, 329, 330, 331, 332, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 352, 353, 354, 355, 356, 357, 358, 359, 360, 361, 362, 363, 364, 365, 366, 367, 368, 369, 370, 371, 372, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384, 385, 386, 387, 388, 389, 390, 391, 392, 393, 394, 395, 396, 397, 398, 399, 400, 401, 402, 403, 404, 405, 406, 407, 408, 409, 410, 411, 412, 413, 414, 415, 416, 417, 418, 419, 420, 421, 422, 423, 424, 425, 426, 427, 428, 429, 430, 431, 432, 433, 434, 435, 436, 437, 438, 439, 440, 441, 442, 443, 444, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 460, 461, 462, 463, 464, 465, 466, 467, 468, 469, 470, 471, 472, 473, 474, 475, 476, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505, 506, 507, 508, 509, 510, 511, 512, 513, 514, 515, 516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 529, 530, 531, 532, 533, 534, 535, 536, 537, 538, 539, 540, 541, 542, 543, 544, 545, 546, 547, 548, 549, 550, 551, 552, 553, 554, 555, 556, 557, 558, 559, 560, 561, 562, 563, 564, 565, 566, 567, 568, 569, 570, 571, 572, 573, 574, 575, 576, 577, 578, 579, 580, 581, 582, 583, 584, 585, 586, 587, 588, 589, 590, 591, 592, 593, 594, 595, 596, 597, 598, 599, 600, 601, 602, 603, 604, 605, 606, 607, 608, 609, 610, 611, 612, 613, 614, 615, 616, 617, 618, 619, 620, 621, 622, 623, 624, 625, 626, 627, 628, 629, 630, 631, 632, 633, 634, 635, 636, 637, 638, 639, 640, 641, 642, 643, 644, 645, 646, 647, 648, 649, 650, 651, 652, 653, 654, 655, 656, 657, 658, 659, 660, 661, 662, 663, 664, 665, 666, 667, 668, 669, 670, 671, 672, 673, 674, 675, 676, 677, 678, 679, 680, 681, 682, 683, 684, 685, 686, 687, 688, 689, 690, 691, 692, 693, 694, 695, 696, 697, 698, 699, 700, 701, 702, 703, 704, 705, 706, 707, 708, 709, 710, 711, 712, 713, 714, 715, 716, 717, 718, 719, 720, 721, 722, 723, 724, 725, 726, 727, 728, 729, 730, 731, 732, 733, 734, 735, 736, 737};

localparam int D_values[638] = {
5, 5, 9, 5, 5, 5, 5, 10, 6, 4, 10, 3, 3, 8, 3, 3, 7, 9, 6, 1, 10, 5, 5, 5, 8, 5, 1, 9, 5, 3, 9, 6, 5, 3, 1, 10, 5, 9, 4, 5, 10, 3, 5, 10, 5, 4, 9, 5, 10, 5, 6, 8, 10, 4, 5, 6, 5, 9, 5, 10, 5, 10, 5, 7, 5, 9, 5, 3, 7, 2, 7, 8, 10, 5, 4, 3, 2, 1, 5, 5, 8, 9, 1, 5, 10, 4, 10, 7, 5, 7, 10, 5, 2, 1, 5, 2, 1, 5, 2, 1, 5, 7, 10, 5, 10, 5, 7, 8, 8, 9, 5, 8, 8, 3, 8, 7, 1, 5, 4, 7, 6, 9, 3, 5, 4, 10, 3, 5, 4, 7, 10, 7, 6, 4, 6, 8, 1, 5, 1, 7, 7, 7, 4, 6, 5, 1, 5, 8, 7, 3, 10, 5, 9, 7, 3, 1, 5, 6, 9, 8, 1, 5, 10, 1, 9, 6, 9, 9, 7, 9, 5, 10, 3, 9, 10, 7, 8, 1, 8, 2, 9, 9, 5, 10, 10, 5, 4, 9, 9, 5, 6, 5, 2, 8, 5, 9, 10, 4, 5, 2, 8, 5, 9, 9, 9, 5, 9, 9, 10, 7, 4, 1, 5, 9, 9, 8, 6, 2, 6, 7, 5, 9, 2, 6, 7, 9, 9, 10, 5, 1, 8, 3, 1, 10, 5, 10, 5, 5, 9, 5, 10, 1, 10, 5, 9, 6, 5, 1, 7, 7, 7, 7, 9, 7, 1, 10, 7, 1, 10, 7, 7, 7, 7, 10, 10, 4, 5, 9, 7, 7, 10, 10, 4, 2, 9, 1, 3, 7, 7, 9, 8, 8, 10, 6, 7, 10, 10, 9, 5, 8, 10, 7, 5, 3, 10, 6, 7, 3, 10, 5, 5, 2, 4, 1, 4, 2, 7, 10, 9, 9, 7, 10, 9, 5, 5, 8, 9, 8, 8, 5, 7, 1, 3, 7, 5, 1, 7, 9, 3, 7, 5, 1, 4, 2, 7, 10, 5, 7, 3, 10, 8, 3, 1, 7, 2, 7, 10, 6, 5, 8, 6, 1, 10, 2, 4, 10, 6, 5, 10, 6, 5, 8, 6, 1, 4, 9, 10, 10, 8, 3, 7, 9, 1, 5, 5, 6, 1, 4, 9, 3, 9, 1, 10, 2, 7, 10, 8, 3, 9, 4, 10, 6, 8, 8, 6, 1, 9, 9, 8, 6, 1, 9, 9, 8, 6, 1, 9, 9, 8, 6, 1, 9, 5, 2, 7, 10, 9, 10, 2, 3, 8, 1, 4, 9, 8, 6, 1, 9, 5, 5, 5, 7, 6, 8, 10, 9, 3, 6, 1, 5, 5, 7, 4, 10, 8, 10, 2, 3, 8, 1, 9, 7, 5, 9, 10, 7, 3, 1, 4, 5, 5, 9, 10, 8, 10, 9, 8, 6, 1, 6, 3, 2, 7, 9, 1, 9, 5, 7, 4, 10, 9, 7, 5, 10, 7, 10, 9, 8, 5, 4, 7, 10, 9, 8, 6, 1, 6, 3, 2, 3, 6, 1, 6, 3, 2, 3, 6, 1, 6, 3, 8, 9, 10, 9, 4, 7, 7, 4, 10, 8, 9, 8, 9, 7, 8, 1, 6, 3, 2, 3, 6, 10, 7, 10, 9, 8, 9, 10, 9, 4, 5, 9, 5, 4, 10, 11, 9, 8, 2, 3, 6, 9, 8, 7, 9, 7, 7, 10, 1, 5, 3, 2, 8, 5, 10, 9, 4, 5, 7, 7, 8, 1, 6, 3, 3, 9, 8, 2, 3, 5, 10, 11, 9, 8, 2, 3, 5, 10, 10, 4, 8, 2, 3, 5, 5, 9, 4, 5, 2, 3, 6, 3, 9, 4, 5, 9, 3, 6, 10, 8, 4, 5, 7, 1, 8, 4, 5, 2, 3, 5, 10, 10, 9, 3, 9, 8, 4, 10, 1, 6, 10, 9, 7, 7, 7, 9, 8, 4};

localparam real M_values[638] = {
64.0, 64.0, 115.0, 64.0, 64.0, 64.0, 64.0, 127.625, 76.625, 51.125, 127.875, 38.375, 38.375, 102.375, 38.375, 38.375, 89.5, 115.0, 76.625, 12.75, 127.375, 64.0, 64.0, 64.0, 102.375, 63.875, 12.75, 114.5, 64.0, 38.375, 114.875, 76.375, 64.0, 38.375, 12.75, 127.125, 64.0, 114.875, 50.875, 64.0, 127.625, 38.125, 64.0, 127.375, 64.0, 51.125, 114.5, 64.0, 127.375, 64.0, 76.625, 101.625, 127.875, 50.875, 64.0, 76.375, 64.0, 114.625, 64.0, 127.375, 64.0, 127.375, 64.0, 89.125, 64.0, 114.5, 64.0, 38.125, 89.5, 25.375, 89.375, 101.375, 127.375, 64.0, 50.875, 38.375, 25.375, 12.75, 64.0, 63.625, 102.375, 114.125, 12.75, 64.0, 127.125, 51.125, 126.625, 89.125, 64.0, 88.75, 127.375, 64.0, 25.375, 12.75, 64.0, 25.375, 12.75, 64.0, 25.375, 12.75, 64.0, 88.75, 127.375, 64.0, 126.625, 63.625, 89.5, 101.125, 101.625, 114.875, 64.0, 101.375, 101.875, 38.375, 101.125, 88.875, 12.75, 64.0, 50.625, 89.0, 76.625, 113.5, 38.0, 63.625, 51.125, 126.125, 38.0, 63.625, 51.125, 88.25, 126.625, 89.0, 76.625, 50.375, 75.875, 101.625, 12.75, 64.0, 12.625, 88.75, 89.125, 89.5, 50.375, 75.875, 63.5, 12.75, 64.0, 100.875, 88.625, 38.125, 127.625, 64.0, 113.5, 88.625, 38.125, 12.75, 64.0, 75.625, 113.875, 101.625, 12.75, 64.0, 125.875, 12.625, 114.125, 76.375, 115.0, 113.0, 88.25, 113.875, 63.5, 127.375, 38.375, 113.125, 126.125, 88.625, 101.625, 12.75, 102.375, 25.125, 113.5, 113.875, 63.5, 127.375, 127.875, 62.75, 50.375, 113.75, 114.125, 63.625, 76.625, 64.0, 25.125, 100.875, 63.25, 114.25, 127.375, 51.125, 62.625, 25.125, 100.875, 63.25, 114.25, 114.625, 115.0, 64.0, 113.0, 113.375, 126.375, 88.75, 50.875, 12.75, 64.0, 112.75, 113.125, 100.875, 75.875, 25.375, 76.375, 89.375, 64.0, 112.75, 25.125, 75.625, 88.5, 114.125, 114.5, 127.625, 64.0, 12.5, 100.375, 37.75, 12.625, 126.625, 63.5, 127.375, 63.875, 64.0, 112.625, 62.75, 125.875, 12.625, 126.625, 63.5, 114.625, 76.625, 64.0, 12.5, 87.75, 88.0, 88.25, 88.5, 114.125, 89.0, 12.75, 127.875, 87.25, 12.5, 125.375, 88.0, 88.25, 88.5, 88.75, 127.125, 127.375, 51.125, 62.25, 112.375, 87.625, 87.875, 125.875, 126.125, 50.625, 25.375, 114.5, 12.75, 38.375, 87.125, 87.375, 112.625, 100.375, 100.625, 126.125, 75.875, 88.75, 127.125, 127.375, 115.0, 64.0, 99.625, 124.875, 87.625, 62.75, 37.75, 126.125, 75.875, 88.75, 38.125, 127.375, 63.875, 64.0, 24.875, 49.875, 12.5, 50.125, 25.125, 88.125, 126.125, 113.875, 114.125, 89.0, 127.375, 115.0, 64.0, 62.125, 99.625, 112.375, 100.125, 100.375, 62.875, 88.25, 12.625, 38.0, 88.875, 63.625, 12.75, 89.5, 111.5, 37.25, 87.125, 62.375, 12.5, 50.125, 25.125, 88.125, 126.125, 63.25, 88.75, 38.125, 127.375, 102.125, 38.375, 12.375, 86.875, 24.875, 87.25, 124.875, 75.125, 62.75, 100.625, 75.625, 12.625, 126.625, 25.375, 50.875, 127.375, 76.625, 64.0, 123.625, 74.375, 62.125, 99.625, 74.875, 12.5, 50.125, 113.0, 125.875, 126.125, 101.125, 38.0, 88.875, 114.5, 12.75, 63.875, 64.0, 74.125, 12.375, 49.625, 111.875, 37.375, 112.375, 12.5, 125.375, 25.125, 88.125, 126.125, 101.125, 38.0, 114.25, 50.875, 127.375, 76.625, 102.375, 98.625, 74.125, 12.375, 111.625, 111.875, 99.625, 74.875, 12.5, 112.75, 113.0, 100.625, 75.625, 12.625, 113.875, 114.125, 101.625, 76.375, 12.75, 115.0, 64.0, 24.625, 86.375, 123.625, 111.5, 124.125, 24.875, 37.375, 99.875, 12.5, 50.125, 113.0, 100.625, 75.625, 12.625, 113.875, 63.375, 63.5, 63.625, 85.5, 76.625, 102.375, 122.875, 110.75, 37.0, 74.125, 12.375, 62.0, 62.125, 87.125, 49.875, 124.875, 100.125, 125.375, 25.125, 37.75, 100.875, 12.625, 113.875, 88.75, 63.5, 114.5, 127.375, 89.375, 38.375, 12.25, 49.125, 61.5, 61.625, 111.125, 123.625, 99.125, 124.125, 111.875, 99.625, 74.875, 12.5, 75.125, 37.625, 25.125, 88.125, 113.5, 12.625, 113.875, 63.375, 88.875, 50.875, 127.375, 114.875, 89.5, 64.0, 116.625, 85.875, 122.875, 110.75, 98.625, 61.75, 47.125, 86.75, 124.125, 111.875, 99.625, 74.875, 12.5, 75.125, 37.625, 25.125, 37.75, 75.625, 12.625, 75.875, 38.0, 25.375, 38.125, 76.375, 12.75, 76.625, 38.375, 97.625, 110.0, 122.375, 110.375, 49.125, 86.125, 86.25, 49.375, 123.625, 94.125, 111.625, 99.375, 112.0, 87.25, 99.875, 12.5, 75.125, 37.625, 25.125, 37.75, 75.625, 119.875, 88.5, 126.625, 114.125, 101.625, 114.5, 127.375, 114.875, 51.125, 64.0, 109.625, 61.0, 48.875, 122.375, 127.75, 110.5, 98.375, 24.625, 37.0, 74.125, 105.5, 99.125, 86.875, 111.875, 87.125, 87.25, 124.875, 12.5, 62.625, 37.625, 25.125, 100.625, 63.0, 126.125, 113.75, 50.625, 63.375, 88.875, 89.0, 101.875, 12.75, 76.625, 38.375, 34.375, 109.375, 97.375, 24.375, 36.625, 61.125, 122.375, 127.375, 110.5, 98.375, 24.625, 37.0, 61.75, 123.625, 123.875, 49.625, 99.375, 24.875, 37.375, 62.375, 59.0, 112.625, 50.125, 62.75, 25.125, 37.75, 75.625, 35.75, 113.75, 50.625, 63.375, 114.25, 38.125, 76.375, 120.375, 102.125, 51.125, 64.0, 84.75, 12.125, 97.125, 48.625, 60.875, 24.375, 36.625, 61.125, 122.375, 115.375, 110.5, 36.875, 110.75, 98.625, 49.375, 123.625, 12.375, 74.375, 124.125, 111.875, 87.125, 87.25, 87.375, 105.875, 100.125, 50.125};

localparam real O_values[638] = {
16.0, 15.875, 15.625, 15.5, 15.375, 15.25, 15.125, 14.875, 14.75, 14.625, 14.5, 14.375, 14.25, 14.125, 14.0, 13.875, 13.75, 13.625, 13.5, 13.375, 13.25, 13.25, 13.125, 13.0, 12.875, 12.75, 12.625, 12.5, 12.5, 12.375, 12.25, 12.125, 12.125, 12.0, 11.875, 11.75, 11.75, 11.625, 11.5, 11.5, 11.375, 11.25, 11.25, 11.125, 11.125, 11.0, 10.875, 10.875, 10.75, 10.75, 10.625, 10.5, 10.5, 10.375, 10.375, 10.25, 10.25, 10.125, 10.125, 10.0, 10.0, 9.875, 9.875, 9.75, 9.75, 9.625, 9.625, 9.5, 9.5, 9.375, 9.375, 9.25, 9.25, 9.25, 9.125, 9.125, 9.0, 9.0, 9.0, 8.875, 8.875, 8.75, 8.75, 8.75, 8.625, 8.625, 8.5, 8.5, 8.5, 8.375, 8.375, 8.375, 8.25, 8.25, 8.25, 8.125, 8.125, 8.125, 8.0, 8.0, 8.0, 7.875, 7.875, 7.875, 7.75, 7.75, 7.75, 7.625, 7.625, 7.625, 7.625, 7.5, 7.5, 7.5, 7.375, 7.375, 7.375, 7.375, 7.25, 7.25, 7.25, 7.125, 7.125, 7.125, 7.125, 7.0, 7.0, 7.0, 7.0, 6.875, 6.875, 6.875, 6.875, 6.75, 6.75, 6.75, 6.75, 6.75, 6.625, 6.625, 6.625, 6.625, 6.5, 6.5, 6.5, 6.5, 6.5, 6.375, 6.375, 6.375, 6.375, 6.375, 6.25, 6.25, 6.25, 6.25, 6.25, 6.125, 6.125, 6.125, 6.125, 6.125, 6.0, 6.0, 6.0, 6.0, 6.0, 5.875, 5.875, 5.875, 5.875, 5.875, 5.875, 5.75, 5.75, 5.75, 5.75, 5.75, 5.75, 5.625, 5.625, 5.625, 5.625, 5.625, 5.625, 5.5, 5.5, 5.5, 5.5, 5.5, 5.5, 5.5, 5.375, 5.375, 5.375, 5.375, 5.375, 5.375, 5.25, 5.25, 5.25, 5.25, 5.25, 5.25, 5.25, 5.25, 5.125, 5.125, 5.125, 5.125, 5.125, 5.125, 5.125, 5.0, 5.0, 5.0, 5.0, 5.0, 5.0, 5.0, 5.0, 4.875, 4.875, 4.875, 4.875, 4.875, 4.875, 4.875, 4.875, 4.75, 4.75, 4.75, 4.75, 4.75, 4.75, 4.75, 4.75, 4.75, 4.625, 4.625, 4.625, 4.625, 4.625, 4.625, 4.625, 4.625, 4.625, 4.5, 4.5, 4.5, 4.5, 4.5, 4.5, 4.5, 4.5, 4.5, 4.375, 4.375, 4.375, 4.375, 4.375, 4.375, 4.375, 4.375, 4.375, 4.375, 4.25, 4.25, 4.25, 4.25, 4.25, 4.25, 4.25, 4.25, 4.25, 4.25, 4.25, 4.125, 4.125, 4.125, 4.125, 4.125, 4.125, 4.125, 4.125, 4.125, 4.125, 4.125, 4.125, 4.0, 4.0, 4.0, 4.0, 4.0, 4.0, 4.0, 4.0, 4.0, 4.0, 4.0, 4.0, 3.875, 3.875, 3.875, 3.875, 3.875, 3.875, 3.875, 3.875, 3.875, 3.875, 3.875, 3.875, 3.875, 3.75, 3.75, 3.75, 3.75, 3.75, 3.75, 3.75, 3.75, 3.75, 3.75, 3.75, 3.75, 3.75, 3.625, 3.625, 3.625, 3.625, 3.625, 3.625, 3.625, 3.625, 3.625, 3.625, 3.625, 3.625, 3.625, 3.625, 3.625, 3.5, 3.5, 3.5, 3.5, 3.5, 3.5, 3.5, 3.5, 3.5, 3.5, 3.5, 3.5, 3.5, 3.5, 3.5, 3.5, 3.375, 3.375, 3.375, 3.375, 3.375, 3.375, 3.375, 3.375, 3.375, 3.375, 3.375, 3.375, 3.375, 3.375, 3.375, 3.375, 3.375, 3.25, 3.25, 3.25, 3.25, 3.25, 3.25, 3.25, 3.25, 3.25, 3.25, 3.25, 3.25, 3.25, 3.25, 3.25, 3.25, 3.25, 3.25, 3.125, 3.125, 3.125, 3.125, 3.125, 3.125, 3.125, 3.125, 3.125, 3.125, 3.125, 3.125, 3.125, 3.125, 3.125, 3.125, 3.125, 3.125, 3.125, 3.125, 3.0, 3.0, 3.0, 3.0, 3.0, 3.0, 3.0, 3.0, 3.0, 3.0, 3.0, 3.0, 3.0, 3.0, 3.0, 3.0, 3.0, 3.0, 2.875, 3.0, 3.0, 2.875, 2.875, 2.875, 2.875, 2.875, 2.875, 2.875, 2.875, 2.875, 2.875, 2.875, 2.875, 2.875, 2.875, 2.875, 2.875, 2.875, 2.875, 2.875, 2.875, 2.875, 2.875, 2.875, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.75, 2.5, 2.625, 2.625, 2.625, 2.625, 2.625, 2.5, 2.625, 2.625, 2.625, 2.625, 2.625, 2.625, 2.625, 2.625, 2.625, 2.625, 2.625, 2.625, 2.625, 2.625, 2.625, 2.625, 2.625, 2.625, 2.625, 2.625, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.375, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.375, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.5, 2.375, 2.375, 2.375, 2.375, 2.25, 2.375, 2.375, 2.375, 2.375, 2.375, 2.25, 2.375, 2.375, 2.375, 2.375, 2.375, 2.375, 2.375, 2.375, 2.375, 2.375, 2.375, 2.375, 2.375, 2.375, 2.375, 2.375, 2.375, 2.375, 2.375, 2.375, 2.375, 2.375, 2.125, 2.25, 2.25, 2.25, 2.25, 2.25, 2.25, 2.125, 2.25, 2.25, 2.25, 2.25, 2.25, 2.25, 2.25, 2.25, 2.25, 2.25, 2.25, 2.25, 2.125, 2.25, 2.25, 2.25, 2.25, 2.25, 2.25, 2.125, 2.25, 2.25, 2.25, 2.25, 2.25, 2.25, 2.125, 2.25, 2.25, 2.25, 2.125, 2.125, 2.125, 2.125, 2.125, 2.125, 2.125, 2.125, 2.125, 2.0, 2.125, 2.125, 2.125, 2.125, 2.125, 2.125, 2.125, 2.125, 2.125, 2.125, 2.125, 2.125, 2.125, 2.0, 2.125, 2.125};

`endif // MMCM_LOOKUP_PARAMS_SVH
