// Lookup table generated from CSV
`ifndef MMCM_LOOKUP_PARAMS_SVH
`define MMCM_LOOKUP_PARAMS_SVH

localparam int desired_freqs[638] = {
100, 101, 102, 103, 104, 105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 214, 215, 216, 217, 218, 219, 220, 221, 222, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 250, 251, 252, 253, 254, 255, 256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 286, 287, 288, 289, 290, 291, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318, 319, 320, 321, 322, 323, 324, 325, 326, 327, 328, 329, 330, 331, 332, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 352, 353, 354, 355, 356, 357, 358, 359, 360, 361, 362, 363, 364, 365, 366, 367, 368, 369, 370, 371, 372, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384, 385, 386, 387, 388, 389, 390, 391, 392, 393, 394, 395, 396, 397, 398, 399, 400, 401, 402, 403, 404, 405, 406, 407, 408, 409, 410, 411, 412, 413, 414, 415, 416, 417, 418, 419, 420, 421, 422, 423, 424, 425, 426, 427, 428, 429, 430, 431, 432, 433, 434, 435, 436, 437, 438, 439, 440, 441, 442, 443, 444, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 460, 461, 462, 463, 464, 465, 466, 467, 468, 469, 470, 471, 472, 473, 474, 475, 476, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 502, 503, 504, 505, 506, 507, 508, 509, 510, 511, 512, 513, 514, 515, 516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 529, 530, 531, 532, 533, 534, 535, 536, 537, 538, 539, 540, 541, 542, 543, 544, 545, 546, 547, 548, 549, 550, 551, 552, 553, 554, 555, 556, 557, 558, 559, 560, 561, 562, 563, 564, 565, 566, 567, 568, 569, 570, 571, 572, 573, 574, 575, 576, 577, 578, 579, 580, 581, 582, 583, 584, 585, 586, 587, 588, 589, 590, 591, 592, 593, 594, 595, 596, 597, 598, 599, 600, 601, 602, 603, 604, 605, 606, 607, 608, 609, 610, 611, 612, 613, 614, 615, 616, 617, 618, 619, 620, 621, 622, 623, 624, 625, 626, 627, 628, 629, 630, 631, 632, 633, 634, 635, 636, 637, 638, 639, 640, 641, 642, 643, 644, 645, 646, 647, 648, 649, 650, 651, 652, 653, 654, 655, 656, 657, 658, 659, 660, 661, 662, 663, 664, 665, 666, 667, 668, 669, 670, 671, 672, 673, 674, 675, 676, 677, 678, 679, 680, 681, 682, 683, 684, 685, 686, 687, 688, 689, 690, 691, 692, 693, 694, 695, 696, 697, 698, 699, 700, 701, 702, 703, 704, 705, 706, 707, 708, 709, 710, 711, 712, 713, 714, 715, 716, 717, 718, 719, 720, 721, 722, 723, 724, 725, 726, 727, 728, 729, 730, 731, 732, 733, 734, 735, 736, 737};

localparam int D_values[638] = {
1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 3, 3, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 3, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 1, 3, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 3, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 3, 3, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 1, 1, 1, 1, 2, 1, 1, 1, 1, 3, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 3, 1, 3, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 3, 3, 1, 1, 1, 2, 1, 1, 1, 1, 2, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 1, 1, 1, 1, 1, 1, 3, 3, 3, 3, 1, 1, 1, 1, 2, 1, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 4, 2, 1, 1, 1, 1, 2, 1, 1, 1, 3, 3, 1, 1, 1, 1, 1, 1, 1, 2, 1, 1, 1, 1, 1, 1, 3, 1, 1, 1, 1, 1, 1, 2, 1, 1, 1, 1, 2, 2, 3, 5, 1, 5, 3, 2, 2, 1, 1, 1, 1, 2, 1, 1, 1, 1, 1, 2, 3, 1, 1, 2, 2, 1, 1, 2, 1, 1, 1, 1, 1, 3, 1, 3, 3, 1, 1, 2, 2, 1, 1, 1, 1, 2, 4, 2, 1, 2, 1, 1, 2, 1, 1, 1, 2, 2, 2, 2, 2, 1, 3, 1, 3, 4, 5, 5, 4, 3, 1, 3, 1, 2, 2, 2, 2, 2, 1, 1, 3, 2, 1, 1, 2, 1, 2, 4, 4, 4, 1, 2, 1, 2, 2, 3, 1, 3, 5, 1, 3, 1, 2, 3, 1, 1, 2, 1, 1, 3, 4, 1, 3, 3, 4, 1, 1, 4, 2, 2, 3, 1, 1, 4, 3, 2, 2, 3, 6, 1, 6, 3, 2, 2, 3, 4, 1, 1, 3, 2, 2, 4, 1, 1, 4, 3, 3, 3, 4, 4, 1, 1, 2, 3, 5, 3, 3, 1, 5, 3, 5, 3, 1, 3, 2, 2, 1, 2, 1, 4, 4, 5, 2, 1, 2, 1, 1, 2, 3, 5, 2, 2, 3, 3, 2, 5, 4, 3, 1, 3, 4, 5, 5, 4, 3, 1, 3, 4, 5, 2, 3, 3, 2, 2, 5, 3, 2, 1, 4, 2, 1, 2, 5, 4, 4, 1, 5, 1, 5, 2, 3, 2, 3, 5, 6, 7, 5, 3, 3, 5, 4, 7, 1, 3, 4, 5, 3, 3, 5, 9, 5, 3};

localparam real M_values[638] = {
6.5, 6.875, 6.625, 6.5, 6.75, 6.5, 6.875, 6.625, 7.125, 6.75, 6.5, 6.875, 6.5, 7.0, 6.5, 7.0, 6.5, 7.125, 6.5, 7.25, 8.625, 7.125, 9.375, 6.875, 12.5, 6.5, 12.75, 7.125, 9.875, 7.625, 6.5, 8.0, 6.875, 8.125, 7.375, 6.625, 7.625, 7.125, 6.625, 7.375, 7.0, 6.625, 7.25, 6.875, 6.625, 7.25, 7.0, 6.625, 7.25, 7.0, 6.75, 6.5, 7.0, 6.875, 6.625, 6.5, 10.125, 6.75, 7.75, 7.0, 6.875, 7.25, 7.125, 7.0, 7.375, 7.25, 7.625, 12.375, 9.25, 8.625, 6.625, 6.5, 6.875, 6.75, 7.125, 7.0, 7.75, 7.25, 7.125, 6.625, 7.375, 6.875, 8.0, 7.5, 6.625, 8.5, 6.875, 19.625, 19.75, 7.0, 8.75, 6.5, 7.875, 6.75, 7.375, 6.625, 7.25, 6.5, 7.125, 8.75, 7.0, 6.625, 6.875, 6.5, 7.75, 7.375, 7.0, 6.625, 15.375, 9.625, 9.25, 6.75, 7.0, 7.25, 8.125, 6.875, 7.125, 7.375, 7.625, 20.375, 9.25, 6.625, 6.875, 8.25, 6.5, 6.75, 7.0, 8.625, 7.75, 6.875, 7.125, 7.625, 6.5, 6.75, 7.25, 7.75, 8.5, 6.875, 7.375, 8.125, 8.875, 6.75, 7.5, 8.5, 10.0, 11.75, 7.375, 9.625, 13.875, 25.375, 6.5, 25.625, 14.125, 9.875, 7.625, 6.625, 10.5, 9.0, 8.0, 7.25, 6.5, 8.875, 8.125, 7.625, 7.125, 6.625, 8.25, 7.75, 7.5, 7.0, 6.75, 6.5, 9.25, 7.375, 7.125, 6.875, 6.625, 7.75, 7.5, 7.25, 7.0, 19.375, 9.875, 9.625, 9.375, 7.125, 10.875, 7.75, 6.625, 8.375, 7.25, 13.375, 21.625, 8.5, 10.0, 7.375, 8.875, 7.125, 7.75, 6.875, 7.5, 6.625, 7.25, 7.875, 9.125, 7.625, 8.875, 6.75, 8.625, 10.5, 7.125, 11.5, 27.125, 27.25, 11.625, 7.25, 10.75, 8.875, 7.0, 9.25, 8.0, 9.625, 8.375, 7.75, 7.125, 6.5, 7.5, 8.5, 7.875, 9.875, 8.25, 11.25, 9.625, 24.625, 15.375, 7.375, 9.75, 7.75, 9.125, 12.875, 8.5, 7.5, 6.5, 12.0, 23.75, 7.25, 9.0, 9.375, 8.0, 8.375, 7.0, 7.375, 9.5, 12.0, 8.5, 8.875, 9.25, 7.5, 7.875, 11.125, 9.0, 6.5, 6.875, 7.625, 8.375, 9.125, 10.25, 11.375, 6.625, 7.75, 8.875, 11.125, 14.875, 20.875, 38.125, 6.75, 38.375, 21.125, 15.125, 11.375, 9.125, 8.0, 6.875, 11.875, 10.75, 9.625, 8.875, 8.125, 7.375, 7.0, 9.75, 12.125, 8.625, 8.25, 10.25, 9.875, 7.125, 6.75, 10.75, 8.375, 8.0, 9.625, 9.25, 7.25, 10.5, 8.5, 28.0, 20.75, 7.75, 9.0, 10.25, 15.625, 7.0, 9.5, 6.625, 9.125, 19.125, 33.375, 12.125, 7.125, 10.5, 8.0, 6.75, 11.0, 9.75, 8.5, 9.375, 10.25, 11.125, 18.875, 10.75, 12.5, 9.5, 12.125, 7.375, 10.0, 31.375, 38.0, 38.125, 31.625, 10.125, 7.5, 12.375, 9.75, 16.875, 11.125, 19.625, 11.625, 10.75, 9.875, 9.0, 10.375, 11.75, 7.25, 8.625, 11.375, 7.75, 14.625, 36.625, 21.125, 10.125, 7.375, 10.625, 7.875, 17.625, 11.625, 10.25, 8.875, 23.875, 32.375, 9.875, 12.25, 8.5, 10.875, 11.375, 9.5, 10.0, 18.125, 8.125, 8.625, 12.0, 12.5, 10.125, 10.625, 26.125, 12.125, 8.75, 9.25, 10.25, 11.25, 12.25, 20.625, 7.875, 8.875, 10.375, 11.875, 15.875, 19.875, 28.375, 52.375, 8.0, 52.625, 28.625, 20.125, 16.125, 12.125, 10.625, 9.125, 8.125, 21.375, 12.75, 11.75, 10.75, 9.75, 9.25, 21.625, 27.875, 11.375, 10.875, 23.875, 22.875, 9.375, 8.875, 19.875, 11.0, 10.5, 12.625, 12.125, 9.5, 31.75, 11.125, 36.625, 27.125, 10.125, 11.75, 17.125, 20.375, 9.125, 12.375, 8.625, 11.875, 24.875, 43.375, 17.375, 9.25, 19.625, 10.375, 8.75, 18.625, 12.625, 11.0, 12.125, 19.875, 22.125, 24.375, 18.875, 21.125, 12.25, 30.125, 9.5, 26.875, 40.375, 47.75, 47.875, 40.625, 27.125, 9.625, 30.625, 12.5, 21.625, 19.375, 25.125, 22.875, 20.625, 12.625, 11.5, 29.375, 19.625, 9.25, 11.0, 20.875, 9.875, 18.625, 46.625, 37.375, 42.125, 9.375, 21.125, 10.0, 22.375, 18.875, 28.375, 11.25, 30.25, 50.5, 12.5, 35.75, 10.75, 25.125, 28.75, 12.0, 12.625, 22.875, 10.25, 10.875, 38.125, 43.625, 12.75, 31.0, 32.875, 46.375, 11.0, 11.625, 44.125, 20.875, 23.375, 35.125, 9.875, 11.125, 39.625, 29.75, 19.875, 24.875, 35.5, 63.625, 10.0, 63.875, 35.75, 25.125, 20.125, 30.25, 40.375, 11.375, 10.125, 36.125, 24.125, 21.625, 45.875, 12.125, 11.5, 48.625, 34.625, 32.75, 30.875, 46.375, 43.875, 11.625, 11.0, 24.625, 37.0, 52.0, 31.25, 33.25, 11.75, 58.875, 35.375, 55.75, 33.5, 12.5, 31.625, 21.125, 25.125, 11.25, 23.875, 10.625, 47.875, 42.625, 53.375, 21.375, 11.375, 24.125, 12.75, 10.75, 22.875, 34.375, 54.0, 21.625, 24.375, 36.625, 34.625, 23.125, 57.875, 46.375, 36.875, 11.625, 32.875, 49.375, 58.375, 58.5, 49.625, 33.125, 11.75, 37.375, 47.125, 59.0, 23.625, 35.5, 37.625, 25.125, 22.375, 56.0, 35.75, 23.875, 11.25, 47.875, 25.375, 12.0, 22.625, 56.625, 45.375, 51.125, 11.375, 60.5, 12.125, 57.125, 22.875, 34.375, 24.375, 36.625, 61.125, 69.125, 80.75, 57.75, 36.875, 34.75, 58.0, 49.375, 86.5, 12.375, 35.0, 49.625, 62.125, 35.125, 37.375, 62.375, 105.875, 58.875, 35.375};

localparam real O_values[638] = {
8.125, 8.5, 8.125, 7.875, 8.125, 7.75, 8.125, 7.75, 8.25, 7.75, 7.375, 7.75, 7.25, 7.75, 7.125, 7.625, 7.0, 7.625, 6.875, 7.625, 9.0, 7.375, 9.625, 7.0, 12.625, 6.5, 12.625, 7.0, 9.625, 7.375, 6.25, 7.625, 6.5, 7.625, 6.875, 6.125, 7.0, 6.5, 6.0, 6.625, 6.25, 5.875, 6.375, 6.0, 5.75, 6.25, 6.0, 5.625, 6.125, 5.875, 5.625, 5.375, 5.75, 5.625, 5.375, 5.25, 8.125, 5.375, 6.125, 5.5, 5.375, 5.625, 5.5, 5.375, 5.625, 5.5, 5.75, 9.25, 6.875, 6.375, 4.875, 4.75, 5.0, 4.875, 5.125, 5.0, 5.5, 5.125, 5.0, 4.625, 5.125, 4.75, 5.5, 5.125, 4.5, 5.75, 4.625, 4.375, 4.375, 4.625, 5.75, 4.25, 5.125, 4.375, 4.75, 4.25, 4.625, 4.125, 4.5, 5.5, 4.375, 4.125, 4.25, 4.0, 4.75, 4.5, 4.25, 4.0, 4.625, 5.75, 5.5, 4.0, 4.125, 4.25, 4.75, 4.0, 4.125, 4.25, 4.375, 3.875, 5.25, 3.75, 3.875, 4.625, 3.625, 3.75, 3.875, 4.75, 4.25, 3.75, 3.875, 4.125, 3.5, 3.625, 3.875, 4.125, 4.5, 3.625, 3.875, 4.25, 4.625, 3.5, 3.875, 4.375, 5.125, 6.0, 3.75, 4.875, 3.5, 6.375, 3.25, 4.25, 3.5, 4.875, 3.75, 3.25, 5.125, 4.375, 3.875, 3.5, 3.125, 4.25, 3.875, 3.625, 3.375, 3.125, 3.875, 3.625, 3.5, 3.25, 3.125, 3.0, 4.25, 3.375, 3.25, 3.125, 3.0, 3.5, 3.375, 3.25, 3.125, 2.875, 4.375, 4.25, 4.125, 3.125, 4.75, 3.375, 2.875, 3.625, 3.125, 2.875, 4.625, 3.625, 4.25, 3.125, 3.75, 3.0, 3.25, 2.875, 3.125, 2.75, 3.0, 3.25, 3.75, 3.125, 3.625, 2.75, 3.5, 4.25, 2.875, 4.625, 3.625, 3.625, 4.625, 2.875, 4.25, 3.5, 2.75, 3.625, 3.125, 3.75, 3.25, 3.0, 2.75, 2.5, 2.875, 3.25, 3.0, 3.75, 3.125, 4.25, 3.625, 4.625, 2.875, 2.75, 3.625, 2.875, 3.375, 2.375, 3.125, 2.75, 2.375, 4.375, 2.875, 2.625, 3.25, 3.375, 2.875, 3.0, 2.5, 2.625, 3.375, 4.25, 3.0, 3.125, 3.25, 2.625, 2.75, 3.875, 3.125, 2.25, 2.375, 2.625, 2.875, 3.125, 3.5, 3.875, 2.25, 2.625, 3.0, 3.75, 2.5, 3.5, 4.25, 2.25, 4.25, 3.5, 2.5, 3.75, 3.0, 2.625, 2.25, 3.875, 3.5, 3.125, 2.875, 2.625, 2.375, 2.25, 3.125, 3.875, 2.75, 2.625, 3.25, 3.125, 2.25, 2.125, 3.375, 2.625, 2.5, 3.0, 2.875, 2.25, 3.25, 2.625, 2.875, 2.125, 2.375, 2.75, 3.125, 2.375, 2.125, 2.875, 2.0, 2.75, 2.875, 2.5, 3.625, 2.125, 3.125, 2.375, 2.0, 3.25, 2.875, 2.5, 2.75, 3.0, 3.25, 2.75, 3.125, 3.625, 2.75, 3.5, 2.125, 2.875, 3.0, 3.625, 3.625, 3.0, 2.875, 2.125, 3.5, 2.75, 2.375, 3.125, 2.75, 3.25, 3.0, 2.75, 2.5, 2.875, 3.25, 2.0, 2.375, 3.125, 2.125, 2.0, 2.5, 2.875, 2.75, 2.0, 2.875, 2.125, 2.375, 3.125, 2.75, 2.375, 2.125, 2.875, 2.625, 3.25, 2.25, 2.875, 3.0, 2.5, 2.625, 2.375, 2.125, 2.25, 3.125, 3.25, 2.625, 2.75, 2.25, 3.125, 2.25, 2.375, 2.625, 2.875, 3.125, 2.625, 2.0, 2.25, 2.625, 3.0, 2.0, 2.5, 2.375, 2.625, 2.0, 2.625, 2.375, 2.5, 2.0, 3.0, 2.625, 2.25, 2.0, 2.625, 3.125, 2.875, 2.625, 2.375, 2.25, 2.625, 2.25, 2.75, 2.625, 2.875, 2.75, 2.25, 2.125, 2.375, 2.625, 2.5, 3.0, 2.875, 2.25, 2.5, 2.625, 2.875, 2.125, 2.375, 2.75, 2.0, 2.375, 2.125, 2.875, 2.0, 2.75, 2.875, 2.5, 2.0, 2.125, 2.25, 2.375, 2.0, 2.125, 2.875, 2.5, 2.75, 2.25, 2.5, 2.75, 2.125, 2.375, 2.75, 2.25, 2.125, 2.0, 2.25, 2.125, 2.125, 2.25, 2.0, 2.125, 2.25, 2.75, 2.375, 2.125, 2.75, 2.5, 2.25, 2.75, 2.5, 2.125, 2.125, 2.0, 2.375, 2.25, 2.125, 2.0, 2.5, 2.0, 2.25, 2.0, 2.25, 2.125, 2.375, 2.0, 2.0, 2.375, 2.125, 2.125, 2.625, 2.5, 2.25, 2.625, 2.0, 2.5, 2.625, 2.375, 2.125, 2.25, 2.625, 2.25, 2.625, 2.125, 2.25, 2.375, 2.25, 2.375, 2.25, 2.125, 2.375, 2.375, 2.0, 2.25, 2.0, 2.0, 2.0, 2.5, 2.375, 2.125, 2.0, 2.125, 2.375, 2.5, 2.0, 2.0, 2.0, 2.25, 2.0, 2.375, 2.375, 2.125, 2.25, 2.375, 2.25, 2.375, 2.25, 2.125, 2.0, 2.25, 2.125, 2.25, 2.125, 2.375, 2.375, 2.0, 2.0, 2.125, 2.25, 2.25, 2.25, 2.125, 2.125, 2.375, 2.0, 2.0, 2.375, 2.125, 2.25, 2.0, 2.25, 2.0, 2.0, 2.0, 2.125, 2.25, 2.375, 2.0, 2.125, 2.125, 2.0, 2.0, 2.25, 2.25, 2.125, 2.125, 2.125, 2.125, 2.25, 2.125, 2.0, 2.25, 2.125, 2.125, 2.25, 2.0, 2.125, 2.25, 2.125, 2.125, 2.125, 2.125, 2.25, 2.25, 2.0, 2.0, 2.125, 2.125, 2.0, 2.125, 2.25, 2.125, 2.0, 2.0, 2.0, 2.25, 2.0, 2.125, 2.125, 2.0, 2.0, 2.0, 2.125, 2.125, 2.125, 2.0, 2.0, 2.0, 2.125, 2.0, 2.0, 2.125, 2.125, 2.125, 2.0, 2.125, 2.125, 2.0, 2.125, 2.125, 2.0, 2.0, 2.0};

`endif // MMCM_LOOKUP_PARAMS_SVH
